module top (
    input wire i_x,
    output wire o_y
);
    assign o_y = i_x;
endmodule