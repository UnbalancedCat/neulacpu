`ifndef MYCPU_VH
    `define MYCPU_VH

    `define BR_BUS_WD       33
    `define FS_TO_DS_BUS_WD 64
    `define DS_TO_ES_BUS_WD 160
    `define ES_TO_MS_BUS_WD 78
    `define MS_TO_WS_BUS_WD 70
    `define WS_TO_RF_BUS_WD 38

    `define DS_TO_FW_BUS_WD 10
    `define ES_TO_FW_BUS_WD 12
    `define MS_TO_FW_BUS_WD 6
    `define FW_TO_ES_BUS_WD 5
    `define MS_TO_ES_BUS_WD 32
    `define WS_TO_ES_BUS_WD 32
`endif
